
module clk_sys (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
